 module top(
input                                sys_clk,
input                                rst_n,
inout                                cmos_scl,         
inout                                cmos_sda,         
input                                cmos_vsync,       
input                                cmos_href,        
input                                cmos_pclk,         
output                               cmos_xclk,         
input [7:0]                          cmos_db,
//ddr                                                           
//output reg                           clk_led               ,
output                               pll_lock               ,
output                               ddr_init_done          ,
output                               ddrphy_rst_done        ,                                                                                                                          
input                                pad_loop_in            ,
input                                pad_loop_in_h          ,
output                               pad_rstn_ch0           ,
output                               pad_ddr_clk_w          ,
output                               pad_ddr_clkn_w         ,
output                               pad_csn_ch0            ,
output [15:0]                        pad_addr_ch0           ,
inout  [16-1:0]                      pad_dq_ch0             ,
inout  [16/8-1:0]                    pad_dqs_ch0            ,
inout  [16/8-1:0]                    pad_dqsn_ch0           ,
output [16/8-1:0]                    pad_dm_rdqs_ch0        ,
output                               pad_cke_ch0            ,
output                               pad_odt_ch0            ,
output                               pad_rasn_ch0           ,
output                               pad_casn_ch0           ,
output                               pad_wen_ch0            ,
output [2:0]                         pad_ba_ch0             ,
output                               pad_loop_out           ,
output                               pad_loop_out_h         ,
//output                               err_flag,   
//hdmi output        
output                             tmds_clk_p,
output                             tmds_clk_n,
output [2:0]                        tmds_data_p,       
output [2:0]                        tmds_data_n,
//caiji output
output  sum_out1 , 
output data_fifo,
input   key,
output cj_clk,
output [7:0]  quotient_1,
output [7:0]  reminder_1,
output   [15:0]  xl_out,


//output xl_out 

output  [4:0]ds_en,
output  [7:0]ds_reg

                       
);

wire [8:0] sum_out1;
wire  caijiclk;
wire  cj_clk;
wire  vs_s;
wire    [8:0 ]data_fifo;
wire    [15:0]  xl_out;
wire  [7:0] sum_out;
wire  [7:0] s_out;
wire [7:0]quotient_1;
wire [7:0]reminder_1;

wire [19:0] d;


wire button_negedge_key3;
wire [3:0] led_eeprom; 
wire[7:0]                       read_data_eep;
parameter MEM_DATA_BITS          = 64;             //external memory user interface data width
parameter ADDR_BITS              = 25;             //external memory user interface address width
parameter BUSRT_BITS             = 10;             //external memory user interface burst width
wire                            wr_burst_data_req;
wire                            wr_burst_finish;
wire                            rd_burst_finish;
wire                            rd_burst_req;
wire                            wr_burst_req;
wire[BUSRT_BITS - 1:0]          rd_burst_len;
wire[BUSRT_BITS - 1:0]          wr_burst_len;
wire[ADDR_BITS - 1:0]           rd_burst_addr;
wire[ADDR_BITS - 1:0]           wr_burst_addr;
wire                            rd_burst_data_valid;
wire[MEM_DATA_BITS - 1 : 0]     rd_burst_data;
wire[MEM_DATA_BITS - 1 : 0]     wr_burst_data;
wire                            read_req;
wire                            read_req_ack;
wire                            read_en;
wire[15:0]                      read_data/*synthesis syn_keep=1*/;
wire                            write_en;
wire[15:0]                      write_data/*synthesis syn_keep=1*/;
wire                            write_req;
wire                            write_req_ack;
wire                            video_clk;         //video pixel clock
wire                            video_clk5x;
wire                            hs;
wire                            vs;
wire                            de;
wire[15:0]                      vout_data;
wire[15:0]                      cmos_16bit_data;
wire                            cmos_16bit_wr;
wire[1:0]                       write_addr_index;
wire[1:0]                       read_addr_index;
wire[9:0]                       lut_index;
wire[31:0]                      lut_data;

wire                            ui_clk;
wire                            ui_clk_sync_rst;
wire                            init_calib_complete;
// Master Write Address
wire [3:0]                      s00_axi_awid;
wire [63:0]                     s00_axi_awaddr;
wire [7:0]                      s00_axi_awlen;    // burst length: 0-255
wire [2:0]                      s00_axi_awsize;   // burst size: fixed 2'b011
wire [1:0]                      s00_axi_awburst;  // burst type: fixed 2'b01(incremental burst)
wire                            s00_axi_awlock;   // lock: fixed 2'b00
wire [3:0]                      s00_axi_awcache;  // cache: fiex 2'b0011
wire [2:0]                      s00_axi_awprot;   // protect: fixed 2'b000
wire [3:0]                      s00_axi_awqos;    // qos: fixed 2'b0000
wire [0:0]                      s00_axi_awuser;   // user: fixed 32'd0
wire                            s00_axi_awvalid;
wire                            s00_axi_awready;
// master write data
wire [63:0]                     s00_axi_wdata;
wire [7:0]                      s00_axi_wstrb;
wire                            s00_axi_wlast;
wire [0:0]                      s00_axi_wuser;
wire                            s00_axi_wvalid;
wire                            s00_axi_wready;
// master write response
wire [3:0]                      s00_axi_bid;
wire [1:0]                      s00_axi_bresp;
wire [0:0]                      s00_axi_buser;
wire                            s00_axi_bvalid;
wire                            s00_axi_bready;
// master read address
wire [3:0]                      s00_axi_arid;
wire [63:0]                     s00_axi_araddr;
wire [7:0]                      s00_axi_arlen;
wire [2:0]                      s00_axi_arsize;
wire [1:0]                      s00_axi_arburst;
wire [1:0]                      s00_axi_arlock;
wire [3:0]                      s00_axi_arcache;
wire [2:0]                      s00_axi_arprot;
wire [3:0]                      s00_axi_arqos;
wire [0:0]                      s00_axi_aruser;
wire                            s00_axi_arvalid;
wire                            s00_axi_arready;
// master read data
wire [3:0]                      s00_axi_rid;
wire [63:0]                     s00_axi_rdata;
wire [1:0]                      s00_axi_rresp;
wire                            s00_axi_rlast;
wire [0:0]                      s00_axi_ruser;
wire                            s00_axi_rvalid;
wire                            s00_axi_rready;
wire                            clk_200MHz;

wire                            hdmi_hs;
wire                            hdmi_vs;
wire                            hdmi_de;
wire[7:0]                       hdmi_r;
wire[7:0]                       hdmi_g;
wire[7:0]                       hdmi_b;
assign  hdmi_hs    = hs;
assign  hdmi_vs     = vs;
assign  hdmi_de    = de;
assign hdmi_r      = {vout_data[15:11],3'd0};
assign hdmi_g      = {vout_data[10:5],2'd0};
assign hdmi_b      = {vout_data[4:0],3'd0};

assign write_en = cmos_16bit_wr;
assign write_data = {cmos_16bit_data[4:0],cmos_16bit_data[10:5],cmos_16bit_data[15:11]};

wire                             sys_clk_g;
wire                             cmos_pclk_g;
wire                             video_clk_w;       
wire                             video_clk5x_w;
wire                             cmos_xclk_w;

wire                             lcd_clk_w;
GTP_CLKBUFG sys_clkbufg
(
  .CLKOUT                    (sys_clk_g                ),
  .CLKIN                     (sys_clk                  )
);
GTP_CLKBUFG cmos_pclkbufg
(
  .CLKOUT                    (cmos_pclk_g              ),
  .CLKIN                     (cmos_pclk                )
);
GTP_CLKBUFG lcd_clkbufg
(
  .CLKOUT                    (lcd_clk                  ),
  .CLKIN                     (lcd_clk_w                )
);
GTP_CLKBUFG cmos_xclkbufg
(
  .CLKOUT                    (cmos_xclk                ),
  .CLKIN                     (cmos_xclk_w              )
);
GTP_CLKBUFG video_clk5xbufg
(
  .CLKOUT                    (video_clk5x               ),
  .CLKIN                     (video_clk5x_w             )
);
GTP_CLKBUFG video_clkbufg
(
  .CLKOUT                    (video_clk                 ),
  .CLKIN                     (video_clk_w               )
);
wire clk_50M;
video_pll video_pll_m0
(
  .clkin1                    (sys_clk_g                ),
  .clkout0                   (video_clk_w              ),
  .clkout1                   (video_clk5x_w            ),
  .clkout2                   (cmos_xclk_w              ),
  .clkout3                   (lcd_clk_w                ),
  .clkout4                   (caiji_clk               ),
  .pll_rst                   (1'b0                     ),
//  .pll_rst                   (~rst_n                     ),
  .pll_lock                  (clk_50M                  )
);

dvi_encoder dvi_encoder_m0
(
	.pixelclk      (video_clk          ),// system clock
	.pixelclk5x    (video_clk5x        ),// system clock x5
	.rstin         (~rst_n             ),// reset
	.blue_din      (hdmi_b            ),// Blue data in
	.green_din     (hdmi_g            ),// Green data in
	.red_din       (hdmi_r            ),// Red data in
	.hsync         (hdmi_hs           ),// hsync data
	.vsync         (hdmi_vs           ),// vsync data
	.de            (hdmi_de         ),// data enable
	.tmds_clk_p    (tmds_clk_p         ),
	.tmds_clk_n    (tmds_clk_n         ),
	.tmds_data_p   (tmds_data_p        ),//rgb
	.tmds_data_n   (tmds_data_n        ) //rgb
);

//I2C master controller
i2c_config i2c_config_m0(
 //.rst                        (~rst_n                   ),
    .rst                        (~ddr_init_done           ),
	.clk                        (sys_clk_g                ),
	.clk_div_cnt                (16'd500                  ),
	.i2c_addr_2byte             (1'b1                     ),
	.lut_index                  (lut_index                ),
	.lut_dev_addr               (lut_data[31:24]          ),
	.lut_reg_addr               (lut_data[23:8]           ),
	.lut_reg_data               (lut_data[7:0]            ),
	.error                      (                         ),
	.done                       (                         ),
	.i2c_scl                    (cmos_scl                 ),
	.i2c_sda                    (cmos_sda                 )
);
//configure look-up table
lut_ov5640_rgb565_1024_768 lut_ov5640_rgb565_1024_768_m0(
	.lut_index                  (lut_index                ),
	.lut_data                   (lut_data                 )
);
//CMOS sensor 8bit data is converted to 16bit data
cmos_8_16bit cmos_8_16bit_m0(
	.rst                        (~rst_n                   ),
	.pclk                       (cmos_pclk_g              ),
	.pdata_i                    (cmos_db                  ),
	.de_i                       (cmos_href                ),
	.pdata_o                    (cmos_16bit_data          ),
	.hblank                     (                         ),
	.de_o                       (cmos_16bit_wr            )
);
//CMOS sensor writes the request and generates the read and write address index
cmos_write_req_gen cmos_write_req_gen_m0(
	.rst                        (~rst_n                   ),
	.pclk                       (cmos_pclk_g              ),
	.cmos_vsync                 (cmos_vsync               ),
	.write_req                  (write_req                ),
	.write_addr_index           (write_addr_index         ),
	.read_addr_index            (read_addr_index          ),
	.write_req_ack              (write_req_ack            )
);

//The video output timing generator and generate a frame read data request
video_timing_data video_timing_data_m0
(
	.video_clk                  (video_clk                ),
	.rst                        (~rst_n                   ),
	.read_req                   (read_req                 ),
	.read_req_ack               (read_req_ack             ),
	.read_en                    (read_en                  ),
	.read_data                  (read_data                ),
	.hs                         (hs                       ),
	.vs                         (vs                       ),
	.de                         (de                       ),
	.vout_data                  (vout_data                )
);
//video frame data read-write control
frame_read_write frame_read_write_m0
(
	.rst                        (~rst_n                   ),
	.mem_clk                    (ui_clk                   ),
	.rd_burst_req               (rd_burst_req             ),
	.rd_burst_len               (rd_burst_len             ),
	.rd_burst_addr              (rd_burst_addr            ),
	.rd_burst_data_valid        (rd_burst_data_valid      ),
	.rd_burst_data              (rd_burst_data            ),
	.rd_burst_finish            (rd_burst_finish          ),
	.read_clk                   (video_clk                ),
	.read_req                   (read_req                 ),
	.read_req_ack               (read_req_ack             ),
	.read_finish                (                         ),
	.read_addr_0                (24'd0                    ), //The first frame address is 0
	.read_addr_1                (24'd2073600              ), //The second frame address is 24'd2073600 ,large enough address space for one frame of video
	.read_addr_2                (24'd4147200              ),
	.read_addr_3                (24'd6220800              ),
	.read_addr_index            (read_addr_index          ),
	.read_len                   (24'd196608               ),//frame size 
	.read_en                    (read_en                  ),
	.read_data                  (read_data                ),

	.wr_burst_req               (wr_burst_req             ),
	.wr_burst_len               (wr_burst_len             ),
	.wr_burst_addr              (wr_burst_addr            ),
	.wr_burst_data_req          (wr_burst_data_req        ),
	.wr_burst_data              (wr_burst_data            ),
	.wr_burst_finish            (wr_burst_finish          ),
	.write_clk                  (cmos_pclk_g              ),
	.write_req                  (write_req                ),
	.write_req_ack              (write_req_ack            ),
	.write_finish               (                         ),
	.write_addr_0               (24'd0                    ),
	.write_addr_1               (24'd2073600              ),
	.write_addr_2               (24'd4147200              ),
	.write_addr_3               (24'd6220800              ),
	.write_addr_index           (write_addr_index         ),
	.write_len                  (24'd196608               ), //frame size  
	.write_en                   (write_en                 ),
	.write_data                 (write_data               )
);
wire                               pll_lock /*synthesis syn_keep=1*/;
wire                               ddr_init_done /*synthesis syn_keep=1*/;
wire                               ddrphy_rst_done /*synthesis syn_keep=1*/;
ddr3 u_ipsl_hmic_h_top (
    .pll_refclk_in        (sys_clk_g      ),
    .top_rst_n         (rst_n          ),   
    .pll_aclk_0           (               ),
    .pll_aclk_1           (ui_clk         ),
    .pll_aclk_2           (               ),
  //  .pll_lock             (      ),
  //  .ddrphy_rst_done      (),
 
  //  .ddrc_init_done       ( ),
  .pll_lock             (pll_lock      ),
    .ddrphy_rst_done      (ddrphy_rst_done),
  //  .ddrphy_rst_done      (ui_clk_sync_rst),
    .ddrc_init_done       (ddr_init_done ),
    .ddrc_rst         (0),    
      
    .areset_1         (0),               
    .aclk_1           (ui_clk),                                                        
    .awid_1           (s00_axi_awid),       
    .awaddr_1         (s00_axi_awaddr),     
    .awlen_1          (s00_axi_awlen),      
    .awsize_1         (s00_axi_awsize),     
    .awburst_1        (s00_axi_awburst),    
    .awlock_1         (s00_axi_awlock),                       
    .awvalid_1        (s00_axi_awvalid),    
    .awready_1        (s00_axi_awready),    
  //  .awurgent_1       (axi_awurgent),  //? 
  //  .awpoison_1       (axi_awpoison),   //?     
    .awurgent_1       (1'b0),  //? 
    .awpoison_1       (1'b0),   //?                 
    .wdata_1          (s00_axi_wdata),      
    .wstrb_1          (s00_axi_wstrb),      
    .wlast_1          (s00_axi_wlast),      
    .wvalid_1         (s00_axi_wvalid),     
    .wready_1         (s00_axi_wready),                       
    .bid_1            (s00_axi_bid),        
    .bresp_1          (s00_axi_bresp),      
    .bvalid_1         (s00_axi_bvalid),     
    .bready_1         (s00_axi_bready),                                    
    .arid_1           (s00_axi_arid     ),  
    .araddr_1         (s00_axi_araddr   ),  
    .arlen_1          (s00_axi_arlen    ),  
    .arsize_1         (s00_axi_arsize   ),  
    .arburst_1        (s00_axi_arburst  ),  
    .arlock_1         (s00_axi_arlock   ),                      
    .arvalid_1        (s00_axi_arvalid  ),  
    .arready_1        (s00_axi_arready  ),  
   // .arpoison_1       (s00_axi_arqos ),   //?   
    .arpoison_1       (1'b0 ),   //?                  
    .rid_1            (s00_axi_rid      ),  
    .rdata_1          (s00_axi_rdata    ),  
    .rresp_1          (s00_axi_rresp    ),  
    .rlast_1          (s00_axi_rlast    ),  
    .rvalid_1         (s00_axi_rvalid   ),  
    .rready_1         (s00_axi_rready   ),  
   // .arurgent_1       (axi_arurgent ),    //?    
    .arurgent_1       (1'b0),    //?        
    .csysreq_1        (1'b1),               
    .csysack_1        (),           
    .cactive_1        (), 
          
    .csysreq_ddrc     (1'b1),
    .csysack_ddrc     (),
    .cactive_ddrc     (),
             
    .pad_loop_in           (pad_loop_in),
    .pad_loop_in_h         (pad_loop_in_h),
    .pad_rstn_ch0          (pad_rstn_ch0),
    .pad_ddr_clk_w         (pad_ddr_clk_w),
    .pad_ddr_clkn_w        (pad_ddr_clkn_w),
    .pad_csn_ch0           (pad_csn_ch0),
    .pad_addr_ch0          (pad_addr_ch0),
    .pad_dq_ch0            (pad_dq_ch0),
    .pad_dqs_ch0           (pad_dqs_ch0),
    .pad_dqsn_ch0          (pad_dqsn_ch0),
    .pad_dm_rdqs_ch0       (pad_dm_rdqs_ch0),
    .pad_cke_ch0           (pad_cke_ch0),
    .pad_odt_ch0           (pad_odt_ch0),
    .pad_rasn_ch0          (pad_rasn_ch0),
    .pad_casn_ch0          (pad_casn_ch0),
    .pad_wen_ch0           (pad_wen_ch0),
    .pad_ba_ch0            (pad_ba_ch0),
    .pad_loop_out          (pad_loop_out),
    .pad_loop_out_h        (pad_loop_out_h)                                
);   
aq_axi_master u_aq_axi_master
	(
      .ARESETN                     (rst_n                                     ),
	 // .ARESETN                     (~ui_clk_sync_rst                          ),
	  .ACLK                        (ui_clk                                    ),
	  .M_AXI_AWID                  (s00_axi_awid                              ),
	  .M_AXI_AWADDR                (s00_axi_awaddr                            ),
	  .M_AXI_AWLEN                 (s00_axi_awlen                             ),
	  .M_AXI_AWSIZE                (s00_axi_awsize                            ),
	  .M_AXI_AWBURST               (s00_axi_awburst                           ),
	  .M_AXI_AWLOCK                (s00_axi_awlock                            ),
	  .M_AXI_AWCACHE               (s00_axi_awcache                           ),
	  .M_AXI_AWPROT                (s00_axi_awprot                            ),
	  .M_AXI_AWQOS                 (s00_axi_awqos                             ),
	  .M_AXI_AWUSER                (s00_axi_awuser                            ),
	  .M_AXI_AWVALID               (s00_axi_awvalid                           ),
	  .M_AXI_AWREADY               (s00_axi_awready                           ),
	  .M_AXI_WDATA                 (s00_axi_wdata                             ),
	  .M_AXI_WSTRB                 (s00_axi_wstrb                             ),
	  .M_AXI_WLAST                 (s00_axi_wlast                             ),
	  .M_AXI_WUSER                 (s00_axi_wuser                             ),
	  .M_AXI_WVALID                (s00_axi_wvalid                            ),
	  .M_AXI_WREADY                (s00_axi_wready                            ),
	  .M_AXI_BID                   (s00_axi_bid                               ),
	  .M_AXI_BRESP                 (s00_axi_bresp                             ),
	  .M_AXI_BUSER                 (s00_axi_buser                             ),
	  .M_AXI_BVALID                (s00_axi_bvalid                            ),
	  .M_AXI_BREADY                (s00_axi_bready                            ),
	  .M_AXI_ARID                  (s00_axi_arid                              ),
	  .M_AXI_ARADDR                (s00_axi_araddr                            ),
	  .M_AXI_ARLEN                 (s00_axi_arlen                             ),
	  .M_AXI_ARSIZE                (s00_axi_arsize                            ),
	  .M_AXI_ARBURST               (s00_axi_arburst                           ),
	  .M_AXI_ARLOCK                (s00_axi_arlock                            ),
	  .M_AXI_ARCACHE               (s00_axi_arcache                           ),
	  .M_AXI_ARPROT                (s00_axi_arprot                            ),
	  .M_AXI_ARQOS                 (s00_axi_arqos                             ),
	  .M_AXI_ARUSER                (s00_axi_aruser                            ),
	  .M_AXI_ARVALID               (s00_axi_arvalid                           ),
	  .M_AXI_ARREADY               (s00_axi_arready                           ),
	  .M_AXI_RID                   (s00_axi_rid                               ),
	  .M_AXI_RDATA                 (s00_axi_rdata                             ),
	  .M_AXI_RRESP                 (s00_axi_rresp                             ),
	  .M_AXI_RLAST                 (s00_axi_rlast                             ),
	  .M_AXI_RUSER                 (s00_axi_ruser                             ),
	  .M_AXI_RVALID                (s00_axi_rvalid                            ),
	  .M_AXI_RREADY                (s00_axi_rready                            ),
	  .MASTER_RST                  (1'b0                                     ),
	  .WR_START                    (wr_burst_req                             ),
	  .WR_ADRS                     ({wr_burst_addr,3'd0}                     ),
	  .WR_LEN                      ({wr_burst_len,3'd0}                      ),
	  .WR_READY                    (                                         ),
	  .WR_FIFO_RE                  (wr_burst_data_req                        ),
	  .WR_FIFO_EMPTY               (1'b0                                     ),
	  .WR_FIFO_AEMPTY              (1'b0                                     ),
	  .WR_FIFO_DATA                (wr_burst_data                            ),
	  .WR_DONE                     (wr_burst_finish                          ),
	  .RD_START                    (rd_burst_req                             ),
	  .RD_ADRS                     ({rd_burst_addr,3'd0}                     ),
	  .RD_LEN                      ({rd_burst_len,3'd0}                      ),
	  .RD_READY                    (                                         ),
	  .RD_FIFO_WE                  (rd_burst_data_valid                      ),
	  .RD_FIFO_FULL                (1'b0                                     ),
	  .RD_FIFO_AFULL               (1'b0                                     ),
	  .RD_FIFO_DATA                (rd_burst_data                            ),
	  .RD_DONE                     (rd_burst_finish                          ),
	  .DEBUG                       (                                         )
);
caiji caiji_1
(
.clk                               (video_clk                                ),
.vout_data                         (vout_data                                ), 
.rst                               (~rst_n                                   ),
. sum_out                          (sum_out1                                 ),
//.en                              (                                         ),
.key                               (key                                      ),
.vs                                (vs                                       ),
.vs_s                              (vs_s                                     )
 );



/*jiance jiance_1(
.clk                               (video_clk                              ),
.sum_out                           (    sumout1                             ), 
.rst                               (~rst_n                                   ),
.sum                               (   data_fifo                           )
 );     */



cj_clk cj_clk_1(
.clk                               (caiji_clk                                ),
.rst                               (~rst_n                                   ),
.cj_clk_r                          (cj_clk                                   )

   );

fifo_in_out fifo_in_out_1 (
.sys_clk                           (      sys_clk_g                        ),         // ʱ���ź�
.cj_clk                            (cj_clk                                   ),
.rst_n                             (~rst_n                                    ),     // ��λ�ź�
.sum1                              (sumout1                                     ),
.vs_s                              (vs_s                                     ),
.data_fifo                         ( data_fifo                               )
);  

chuli chuli_1(
.clk(sys_clk_g ),
.data(data_fifo  ),
.en( rdreq ),
.rst(~rst_n),
//.xl_out(xl_out),
.sum_out(sum_out),
.s_out(s_out)

   );

/*divider_module divider_module_1 (
.dividend                              ( sum_out                               ),
.divisor                                (s_out                              ),
.clk                                   (caiji_clk                               ),
.rst                                   (rst_n                             ),
.quotient                              (quotient_1                              ),
.reminder                               (reminder_1                           )
);  */


multiple8 multiple8_1(
.clk(   video_clk                                                      ),
.rst_n(~ rst_n                                                         ),
.mul_a(s_out                                                          ),
.mul_b(3'd6                                                          ),
.result( xl_out                                                       )
    );


/*xianshi xianshi_1(
.d(d),
.s_out(s_out)
);*/

assign d[19:16] =  xl_out/100%10;//dis/10000;    // ��λ
assign d[15:12] =  xl_out/10%10;//dis/1000%10;  // ʮλ
assign d[11:8]  = xl_out%10;//dis/100%10;   // ��λ
assign d[7:4]   =  xl_out*10%10;//dis/10%10;    // 0.1
assign d[3:0]   = xl_out*100%10;//dis%10;       // 0.01
   
wire  [4:0]ds_en ;
wire  [7:0]ds_reg ;
translator translator_1(
.clk                               (    sys_clk_g               ),
.res_n                             (     rst_n            ),
.num1                (            d[19:16]                               ),//��λ
.num2                (            d[15:12]                               ), //ʮλ
.num3                (            d[11:8]                                ),//��λ
.num4                (            d[7:4]                                 ), //0.1
.num5                (            d[3:0]                                 ), //0.01
.ds_en               (            ds_en                                   ),//5λ�����ʹ��,�����λѡ��ѡ��ǰҪ��ʾ�������
.ds_reg              (            ds_reg                               )	//����ܶ�ѡ����ǰҪ��ʾ������
);


endmodule